// two multiplexers were not implemented in the supporting modules
// They are ALU operand 2 and writeDestination multiplexer
// TODO Implement them here and connect the wiring properly
module EX_Stage();




endmodule
