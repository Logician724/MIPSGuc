module ALU_Control(aluOp, funct, aluControlInput);

input [:] aluOp;
input [5:0] funct;

output [3:0] aluControlInput;




endmodule
