module EX_Stage();




endmodule
